`ifndef KEI_I2C_CONFIGS_SVH
`define KEI_I2C_CONFIGS_SVH

`include "kei_i2c_defines.svh"
`include "kei_i2c_config.sv"

`endif // KEI_I2C_CONFIGS_SVH
