
`ifndef KEI_I2C_VIRTUAL_SEQUENCES_SVH
`define KEI_I2C_VIRTUAL_SEQUENCES_SVH

`include "kei_i2c_base_virtual_sequence.sv" 
`include "kei_i2c_quick_reg_access_virt_seq.sv" 
`include "kei_i2c_master_directed_interrupt_virt_seq.sv" 
`include "kei_i2c_master_directed_write_packet_virt_seq.sv" 
`include "kei_i2c_master_directed_read_packet_virt_seq.sv" 

`endif // KEI_I2C_VIRTUAL_SEQUENCES_SVH

