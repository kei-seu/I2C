
`ifndef KEI_I2C_USER_ELEMENT_SEQUENCES_SVH
`define KEI_I2C_USER_ELEMENT_SEQUENCES_SVH

`include "kei_apb_write_nocheck_packet_seq.sv"

`include "kei_apb_noread_packet_seq.sv"

`endif // KEI_I2C_USER_ELEMENT_SEQUENCES_SVH

