
`ifndef KEI_I2C_USER_TESTS_SVH
`define KEI_I2C_USER_TESTS_SVH

`include "kei_i2c_master_address_cg_test.sv"

`endif // KEI_I2C_USER_TESTS_SVH

