

`ifndef KEI_I2C_CGM_SV
`define KEI_I2C_CGM_SV

// Coverage Model
class kei_i2c_cgm extends uvm_component;
   
  // TODO
  // Covergroup definition below

  // Analysis import declarion below

  `uvm_component_utils(kei_i2c_cgm)

  function new(string name = "kei_i2c_cgm", uvm_component parent = null);
    super.new(name, parent);
  endfunction

endclass


`endif // KEI_I2C_CGM_SV
