
`ifndef KEI_I2C_USER_ELEMENT_SEQUENCES_SVH
`define KEI_I2C_USER_ELEMENT_SEQUENCES_SVH


`endif // KEI_I2C_USER_ELEMENT_SEQUENCES_SVH

