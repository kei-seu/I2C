
`ifndef KEI_I2C_TESTS_SVH
`define KEI_I2C_TESTS_SVH

`include "kei_i2c_base_test.sv"
`include "kei_i2c_quick_reg_access_test.sv"
`include "kei_i2c_master_directed_interrupt_test.sv"
`include "kei_i2c_master_directed_write_packet_test.sv"
`include "kei_i2c_master_directed_read_packet_test.sv"
`include "kei_i2c_reg_access_test.sv"
`include "kei_i2c_reg_bit_bash_test.sv"
`include "kei_i2c_reg_hw_reset_test.sv"

`endif // KEI_I2C_TESTS_SVH
