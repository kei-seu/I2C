
`ifndef KEI_I2C_ELEMENT_SEQUENCES_SVH
`define KEI_I2C_ELEMENT_SEQUENCES_SVH

`include "kei_apb_base_sequence.sv"
`include "kei_apb_config_seq.sv"
`include "kei_apb_tx_seq.sv"
`include "kei_apb_rx_seq.sv"
`include "kei_apb_wait_empty_seq.sv"
`include "kei_apb_intr_enable_seq.sv"

`include "kei_i2c_slave_base_sequence.sv"
`include "kei_i2c_slave_rx_seq.sv"


`endif // KEI_I2C_ELEMENT_SEQUENCES_SVH
