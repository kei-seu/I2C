
`ifndef KEI_I2C_USER_TESTS_SVH
`define KEI_I2C_USER_TESTS_SVH

`include "kei_i2c_master_address_cg_test.sv"

`include "kei_i2c_master_ss_cnt_test.sv"
`include "kei_i2c_master_fs_cnt_test.sv"
`include "kei_i2c_master_hs_cnt_test.sv"

`endif // KEI_I2C_USER_TESTS_SVH

