
`ifndef KEI_I2C_VIRTUAL_SEQUENCES_SVH
`define KEI_I2C_VIRTUAL_SEQUENCES_SVH

`include "kei_i2c_base_virtual_sequence.sv" 
`include "kei_i2c_quick_reg_access_virt_seq.sv" 
`include "kei_i2c_directed_tx_virt_seq.sv" 
`include "kei_i2c_directed_rx_virt_seq.sv" 

`endif // KEI_I2C_VIRTUAL_SEQUENCES_SVH

