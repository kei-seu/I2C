
`ifndef KEI_I2C_USER_VIRTUAL_SEQUENCES_SVH
`define KEI_I2C_USER_VIRTUAL_SEQUENCES_SVH

`include "kei_i2c_master_address_cg_virt_seq.sv"


`endif // KEI_I2C_USER_VIRTUAL_SEQUENCES_SVH

